library ieee;
use ieee.std_logic_1164.all;
use work.dadda_utils.all;
use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;

entity dadda_multi is
  port(
    a: in std_logic_vector(16 downto 0);
    b: in std_logic_vector(16 downto 0);
    p: out std_logic_vector(33 downto 0)
  );
end dadda_multi;

architecture dadda_multi_arch of dadda_multi is
-- Signals having all the parital products
signal l1: std_logic_vector(16 downto 0);
signal l2: std_logic_vector(16 downto 0);
signal l3: std_logic_vector(16 downto 0);
signal l4: std_logic_vector(16 downto 0);
signal l5: std_logic_vector(16 downto 0);
signal l6: std_logic_vector(16 downto 0);
signal l7: std_logic_vector(16 downto 0);
signal l8: std_logic_vector(16 downto 0);
signal l9: std_logic_vector(16 downto 0);
signal l10: std_logic_vector(16 downto 0);
signal l11: std_logic_vector(16 downto 0);
signal l12: std_logic_vector(16 downto 0);
signal l13: std_logic_vector(16 downto 0);
signal l14: std_logic_vector(16 downto 0);
signal l15: std_logic_vector(16 downto 0);
signal l16: std_logic_vector(16 downto 0);
signal l17: std_logic_vector(16 downto 0);
-- Contains the extra partial products which arise due to change to signed dadda multipler
signal extra_pp: std_logic_vector(1 downto 0); 

--Step 1 in Dadda reduction to 13 wires
signal s1_1: std_logic_vector(32 downto 0);	
signal s1_2: std_logic_vector(31 downto 1);
signal s1_3: std_logic_vector(30 downto 2);
signal s1_4: std_logic_vector(29 downto 3);
signal s1_5: std_logic_vector(28 downto 4);
signal s1_6: std_logic_vector(27 downto 5);
signal s1_7: std_logic_vector(26 downto 6);	
signal s1_8: std_logic_vector(25 downto 7);
signal s1_9: std_logic_vector(24 downto 8);
signal s1_10: std_logic_vector(23 downto 9);
signal s1_11: std_logic_vector(22 downto 10);
signal s1_12: std_logic_vector(21 downto 11);
signal s1_13: std_logic_vector(21 downto 12);


--Step 2 in Dadda reduction to 9 wires
signal s2_1: std_logic_vector(32 downto 0);	
signal s2_2: std_logic_vector(31 downto 1);
signal s2_3: std_logic_vector(30 downto 2);
signal s2_4: std_logic_vector(29 downto 3);
signal s2_5: std_logic_vector(28 downto 4);
signal s2_6: std_logic_vector(27 downto 5);
signal s2_7: std_logic_vector(26 downto 6);	
signal s2_8: std_logic_vector(25 downto 7);
signal s2_9: std_logic_vector(25 downto 8);

--Step 3 in Dadda reduction to 6 wires
signal s3_1: std_logic_vector(32 downto 0);	
signal s3_2: std_logic_vector(31 downto 1);
signal s3_3: std_logic_vector(30 downto 2);
signal s3_4: std_logic_vector(29 downto 3);
signal s3_5: std_logic_vector(28 downto 4);
signal s3_6: std_logic_vector(28 downto 5);

--Step 4 in Dadda reduction to 4 wires
signal s4_1: std_logic_vector(32 downto 0);	
signal s4_2: std_logic_vector(31 downto 1);
signal s4_3: std_logic_vector(30 downto 2);
signal s4_4: std_logic_vector(30 downto 3);

--Step 5 in Dadda reduction to 3 wires
signal s5_1: std_logic_vector(32 downto 0);	
signal s5_2: std_logic_vector(31 downto 1);
signal s5_3: std_logic_vector(31 downto 2);

--Step 6 in Dadda reduction to 2 wires
signal s6_1: std_logic_vector(32 downto 0);	
signal s6_2: std_logic_vector(32 downto 0);

signal a_not : std_logic_vector(15 downto 0);

begin
	a_not(15 downto 0) <= not a(15 downto 0);
	-- Partial products in terms of inputs a and b
	l1(15 downto 0) <= and_16b(b(0),a(15 downto 0));
	l1(16) <= a(16) and (not b(0));
	l2(15 downto 0) <= and_16b(b(1),a(15 downto 0));
	l2(16) <= a(16) and (not b(1));
	l3(15 downto 0) <= and_16b(b(2),a(15 downto 0));
	l3(16) <= a(16) and (not b(2));
	l4(15 downto 0) <= and_16b(b(3),a(15 downto 0));
	l4(16) <= a(16) and (not b(3));
	l5(15 downto 0) <= and_16b(b(4),a(15 downto 0));
	l5(16) <= a(16) and (not b(4));
	l6(15 downto 0) <= and_16b(b(5),a(15 downto 0));
	l6(16) <= a(16) and (not b(5));
	l7(15 downto 0) <= and_16b(b(6),a(15 downto 0));
	l7(16) <= a(16) and (not b(6));
	l8(15 downto 0) <= and_16b(b(7),a(15 downto 0));
	l8(16) <= a(16) and (not b(7));
	l9(15 downto 0) <= and_16b(b(8),a(15 downto 0));
	l9(16) <= a(16) and (not b(8));
	l10(15 downto 0) <= and_16b(b(9),a(15 downto 0));
	l10(16) <= a(16) and (not b(9));
	l11(15 downto 0) <= and_16b(b(10),a(15 downto 0));
	l11(16) <= a(16) and (not b(10));
	l12(15 downto 0) <= and_16b(b(11),a(15 downto 0));
	l12(16) <= a(16) and (not b(11));
	l13(15 downto 0) <= and_16b(b(12),a(15 downto 0));
	l13(16) <= a(16) and (not b(12));
	l14(15 downto 0) <= and_16b(b(13),a(15 downto 0));
	l14(16) <= a(16) and (not b(13));
	l15(15 downto 0) <= and_16b(b(14),a(15 downto 0));
	l15(16) <= a(16) and (not b(14));
	l16(15 downto 0) <= and_16b(b(15),a(15 downto 0));
	l16(16) <= a(16) and (not b(15));
	l17(15 downto 0) <= and_16b(b(16),a_not(15 downto 0));
	l17(16) <= a(16) or b(16);

	extra_pp(0) <= a(16) xor b(16);
	extra_pp(1) <= a(16) and b(16);

	--Step 1 Dadda Reduction 

	--Line 1 in 13 wires after 1st reduction

	s1_1(12 downto 0) <= l1(12 downto 0);
	s1_1(13) <= sum_2b(l1(13),l2(12));
	s1_1(14) <= sum_3b(l1(14),l2(13),l3(12));
	s1_1(15) <= sum_3b(l1(15),l2(14),l3(13));
	s1_1(16) <= sum_3b(extra_pp(0),l1(16),l2(15));
	s1_1(17) <= sum_3b(extra_pp(1),l2(16),l3(15));
	s1_1(18) <= sum_3b(l3(16),l4(15),l5(14));
	s1_1(19) <= sum_3b(l4(16),l5(15),l6(14));
	s1_1(20) <= sum_3b(l5(16),l6(15),l7(14));
	s1_1(21) <= l6(16);
	s1_1(22) <= l7(16);
	s1_1(23) <= l8(16);
	s1_1(24) <= l9(16);
	s1_1(25) <= l10(16);
	s1_1(26) <= l11(16);
	s1_1(27) <= l12(16);
	s1_1(28) <= l13(16);
	s1_1(29) <= l14(16);
	s1_1(30) <= l15(16);
	s1_1(31) <= l16(16);
	s1_1(32) <= l17(16);

	--Line 2 in 13 wires after 1st reduction

	s1_2(12 downto 1) <= l2(11 downto 0);
	s1_2(13) <= l3(11);
	s1_2(14) <= carry_2b(l1(13),l2(12));
	s1_2(15) <= carry_3b(l1(14),l2(13),l3(12));
	s1_2(16) <= carry_3b(l1(15),l2(14),l3(13));
	s1_2(17) <= carry_3b(extra_pp(0),l1(16),l2(15));
	s1_2(18) <= carry_3b(extra_pp(1),l2(16),l3(15));
	s1_2(19) <= carry_3b(l3(16),l4(15),l5(14));
	s1_2(20) <= carry_3b(l4(16),l5(15),l6(14));
	s1_2(21) <= carry_3b(l5(16),l6(15),l7(14));
	s1_2(22) <= l8(15);
	s1_2(23) <= l9(15);
	s1_2(24) <= l10(15);
	s1_2(25) <= l11(15);
	s1_2(26) <= l12(15);
	s1_2(27) <= l13(15);
	s1_2(28) <= l14(15);
	s1_2(29) <= l15(15);
	s1_2(30) <= l16(15);
	s1_2(31) <= l17(15);

	--Line 3 in 13 wires after 1st reduction

	s1_3(12 downto 2) <= l3(10 downto 0);
	s1_3(13) <= l4(10);
	s1_3(14) <= sum_2b(l4(11),l5(10));
	s1_3(15) <= sum_3b(l4(12),l5(11),l6(10));
	s1_3(16) <= sum_3b(l3(14),l4(13),l5(12));
	s1_3(17) <= sum_3b(l4(14),l5(13),l6(12));
	s1_3(18) <= sum_3b(l6(13),l7(12),l8(11));
	s1_3(19) <= sum_3b(l7(13),l8(12),l9(11));
	s1_3(20) <= l8(13);
	s1_3(21) <= l7(15);
	s1_3(22) <= l9(14); 
	s1_3(23) <= l10(14);
	s1_3(24) <= l11(14);
	s1_3(25) <= l12(14);
	s1_3(26) <= l13(14);
	s1_3(27) <= l14(14);
	s1_3(28) <= l15(14);
	s1_3(29) <= l16(14);
	s1_3(30) <= l17(14);

	--Line 4 in 13 wires after 1st reduction

	s1_4(12 downto 3) <= l4(9 downto 0);
	s1_4(13) <= l5(9);
	s1_4(14) <= l6(9);
	s1_4(15) <= carry_2b(l4(11),l5(10));
	s1_4(16) <= carry_3b(l4(12),l5(11),l6(10));
	s1_4(17) <= carry_3b(l3(14),l4(13),l5(12));
	s1_4(18) <= carry_3b(l4(14),l5(13),l6(12));
	s1_4(19) <= carry_3b(l6(13),l7(12),l8(11));
	s1_4(20) <= carry_3b(l7(13),l8(12),l9(11));
	s1_4(21) <= l8(14);
	s1_4(22) <= l10(13); 
	s1_4(23) <= l11(13);
	s1_4(24) <= l12(13);
	s1_4(25) <= l13(13);
	s1_4(26) <= l14(13);
	s1_4(27) <= l15(13);
	s1_4(28) <= l16(13);
	s1_4(29) <= l17(13);

		--Line 5 in 13 wires after 1st reduction

	s1_5(12 downto 4) <= l5(8 downto 0);
	s1_5(13) <= l6(8);
	s1_5(14) <= l7(8);
	s1_5(15) <= sum_2b(l7(9),l8(8));
	s1_5(16) <= sum_3b(l6(11),l7(10),l8(9));
	s1_5(17) <= sum_3b(l7(11),l8(10),l9(9));
	s1_5(18) <= sum_3b(l9(10),l10(9),l11(8));
	s1_5(19) <= l10(10);
	s1_5(20) <= l9(12);
	s1_5(21) <= l9(13);
	s1_5(22) <= l11(12); 
	s1_5(23) <= l12(12);
	s1_5(24) <= l13(12);
	s1_5(25) <= l14(12);
	s1_5(26) <= l15(12);
	s1_5(27) <= l16(12);
	s1_5(28) <= l17(12);


	--Line 6 in 13 wires after 1st reduction

	s1_6(12 downto 5) <= l6(7 downto 0);
	s1_6(13) <= l7(7);
	s1_6(14) <= l8(7);
	s1_6(15) <= l9(7);
	s1_6(16) <= carry_2b(l7(9),l8(8));
	s1_6(17) <= carry_3b(l6(11),l7(10),l8(9));
	s1_6(18) <= carry_3b(l7(11),l8(10),l9(9));
	s1_6(19) <= carry_3b(l9(10),l10(9),l11(8));
	s1_6(20) <= l10(11);
	s1_6(21) <= l10(12);
	s1_6(22) <= l12(11);
	s1_6(23) <= l13(11); 
	s1_6(24) <= l14(11);
	s1_6(25) <= l15(11);
	s1_6(26) <= l16(11);
	s1_6(27) <= l17(11);

	--Line 7 in 13 wires after 1st reduction

	s1_7(12 downto 6) <= l7(6 downto 0);
	s1_7(13) <= l8(6);
	s1_7(14) <= l9(6);
	s1_7(15) <= l10(6);
	s1_7(16) <= sum_3b(l9(8),l10(7),l11(6));
	s1_7(17) <= sum_3b(l10(8),l11(7),l12(6));
	s1_7(18) <= l12(7);
	s1_7(19) <= l11(9);
	s1_7(20) <= l11(10);
	s1_7(21) <= l11(11);
	s1_7(22) <= l13(10);
	s1_7(23) <= l14(10); 
	s1_7(24) <= l15(10);
	s1_7(25) <= l16(10);
	s1_7(26) <= l17(10);


	--Line 8 in 13 wires after 1st reduction

	s1_8(12 downto 7) <= l8(5 downto 0);
	s1_8(13) <= l9(5);
	s1_8(14) <= l10(5);
	s1_8(15) <= l11(5);
	s1_8(16) <= l12(5);
	s1_8(17) <= carry_3b(l9(8),l10(7),l11(6));
	s1_8(18) <= carry_3b(l10(8),l11(7),l12(6));
	s1_8(19) <= l12(8);
	s1_8(20) <= l12(9);
	s1_8(21) <= l12(10);
	s1_8(22) <= l14(9);
	s1_8(23) <= l15(9); 
	s1_8(24) <= l16(9);
	s1_8(25) <= l17(9);	

	--Line 9 in 13 wires after 1st reduction

	s1_9(12 downto 8) <= l9(4 downto 0);
	s1_9(13) <= l10(4);
	s1_9(14) <= l11(4);
	s1_9(15) <= l12(4);
	s1_9(16) <= l13(4);
	s1_9(17) <= l13(5);
	s1_9(18) <= l13(6);
	s1_9(19) <= l13(7);
	s1_9(20) <= l13(8);
	s1_9(21) <= l13(9);
	s1_9(22) <= l15(8);
	s1_9(23) <= l16(8); 
	s1_9(24) <= l17(8);	


	--Line 10 in 13 wires after 1st reduction

	s1_10(12 downto 9) <= l10(3 downto 0);
	s1_10(13) <= l11(3);
	s1_10(14) <= l12(3);
	s1_10(15) <= l13(3);
	s1_10(16) <= l14(3);
	s1_10(17) <= l14(4);
	s1_10(18) <= l14(5);
	s1_10(19) <= l14(6);
	s1_10(20) <= l14(7);
	s1_10(21) <= l14(8);
	s1_10(22) <= l16(7);
	s1_10(23) <= l17(7); 	

	--Line 11 in 13 wires after 1st reduction

	s1_11(12 downto 10) <= l11(2 downto 0);
	s1_11(13) <= l12(2);
	s1_11(14) <= l13(2);
	s1_11(15) <= l14(2);
	s1_11(16) <= l15(2);
	s1_11(17) <= l15(3);
	s1_11(18) <= l15(4);
	s1_11(19) <= l15(5);
	s1_11(20) <= l15(6);
	s1_11(21) <= l15(7);
	s1_11(22) <= l17(6);

	--Line 12 in 13 wires after 1st reduction

	s1_12(12 downto 11) <= l12(1 downto 0);
	s1_12(13) <= l13(1);
	s1_12(14) <= l14(1);
	s1_12(15) <= l15(1);
	s1_12(16) <= l16(1);
	s1_12(17) <= l16(2);
	s1_12(18) <= l16(3);
	s1_12(19) <= l16(4);
	s1_12(20) <= l16(5);
	s1_12(21) <= l16(6);

--Line 13 in 13 wires after 1st reduction

	s1_13(12) <= l13(0);
	s1_13(13) <= l14(0);
	s1_13(14) <= l15(0);
	s1_13(15) <= l15(0);
	s1_13(16) <= l17(0);
	s1_13(17) <= l17(1);
	s1_13(18) <= l17(2);
	s1_13(19) <= l17(3);
	s1_13(20) <= l17(4);
	s1_13(21) <= l17(5);

--Line 1 in 9 wires after 2nd reduction
	s2_1(8 downto 0) <= s1_1(8 downto 0);
	s2_1(9) <= sum_2b(s1_1(9),s1_2(9));
	s2_1(10) <= sum_3b(s1_1(10),s1_2(10),s1_3(10));
	s2_1(11) <= sum_3b(s1_1(11),s1_2(11),s1_3(11));	
	s2_1(12) <= sum_3b(s1_1(12),s1_2(12),s1_3(12));
	s2_1(13) <= sum_3b(s1_1(13),s1_2(13),s1_3(13));
	s2_1(14) <= sum_3b(s1_1(14),s1_2(14),s1_3(14));
	s2_1(15) <= sum_3b(s1_1(15),s1_2(15),s1_3(15));
	s2_1(16) <= sum_3b(s1_1(16),s1_2(16),s1_3(16));
	s2_1(17) <= sum_3b(s1_1(17),s1_2(17),s1_3(17));
	s2_1(18) <= sum_3b(s1_1(18),s1_2(18),s1_3(18));
	s2_1(19) <= sum_3b(s1_1(19),s1_2(19),s1_3(19));
	s2_1(20) <= sum_3b(s1_1(20),s1_2(20),s1_3(20));
	s2_1(21) <= sum_3b(s1_1(21),s1_2(21),s1_3(21));
	s2_1(22) <= sum_3b(s1_1(22),s1_2(22),s1_3(22));
	s2_1(23) <= sum_3b(s1_1(23),s1_2(23),s1_3(23));
	s2_1(24) <= sum_3b(s1_1(24),s1_2(24),s1_3(24));
	s2_1(32 downto 25 ) <= s1_1(32 downto 25);

	--Line 2 in 9 wires after 2nd reduction
	s2_2(8 downto 1) <= s1_2(8 downto 1);
	s2_2(9) <= s1_3(9);
	s2_2(10) <= carry_2b(s1_1(9),s1_2(9));
	s2_2(11) <= carry_3b(s1_1(10),s1_2(10),s1_3(10));
	s2_2(12) <= carry_3b(s1_1(11),s1_2(11),s1_3(11));	
	s2_2(13) <= carry_3b(s1_1(12),s1_2(12),s1_3(12));
	s2_2(14) <= carry_3b(s1_1(13),s1_2(13),s1_3(13));
	s2_2(15) <= carry_3b(s1_1(14),s1_2(14),s1_3(14));
	s2_2(16) <= carry_3b(s1_1(15),s1_2(15),s1_3(15));
	s2_2(17) <= carry_3b(s1_1(16),s1_2(16),s1_3(16));
	s2_2(18) <= carry_3b(s1_1(17),s1_2(17),s1_3(17));
	s2_2(19) <= carry_3b(s1_1(18),s1_2(18),s1_3(18));
	s2_2(20) <= carry_3b(s1_1(19),s1_2(19),s1_3(19));
	s2_2(21) <= carry_3b(s1_1(20),s1_2(20),s1_3(20));
	s2_2(22) <= carry_3b(s1_1(21),s1_2(21),s1_3(21));
	s2_2(23) <= carry_3b(s1_1(22),s1_2(22),s1_3(22));
	s2_2(24) <= carry_3b(s1_1(23),s1_2(23),s1_3(23));
	s2_2(25) <= carry_3b(s1_1(24),s1_2(24),s1_3(24));
	s2_2(31 downto 26 ) <= s1_2(31 downto 26);

	--Line 3 in 9 wires after 2nd reduction
	s2_3(8 downto 2) <= s1_3(8 downto 2);
	s2_3(9) <= s1_4(9);
	s2_3(10) <= sum_2b(s1_4(10),s1_5(10));
	s2_3(11) <= sum_3b(s1_4(11),s1_5(11),s1_6(11));
	s2_3(12) <= sum_3b(s1_4(12),s1_5(12),s1_6(12));
	s2_3(13) <= sum_3b(s1_4(13),s1_5(13),s1_6(13));
	s2_3(14) <= sum_3b(s1_4(14),s1_5(14),s1_6(14));
	s2_3(15) <= sum_3b(s1_4(15),s1_5(15),s1_6(15));
	s2_3(16) <= sum_3b(s1_4(16),s1_5(16),s1_6(16));
	s2_3(17) <= sum_3b(s1_4(17),s1_5(17),s1_6(17));
	s2_3(18) <= sum_3b(s1_4(18),s1_5(18),s1_6(18));
	s2_3(19) <= sum_3b(s1_4(19),s1_5(19),s1_6(19));
	s2_3(20) <= sum_3b(s1_4(20),s1_5(20),s1_6(20));
	s2_3(21) <= sum_3b(s1_4(21),s1_5(21),s1_6(21));
	s2_3(22) <= sum_3b(s1_4(22),s1_5(22),s1_6(22));
	s2_3(23) <= sum_3b(s1_4(23),s1_5(23),s1_6(23));
	s2_3(24) <= s1_4(24);
	s2_3(25) <= s1_2(25);
	s2_3(30 downto 26 ) <= s1_3(30 downto 26);

	--Line 4 in 9 wires after 2nd reduction
	s2_4(8 downto 3) <= s1_4(8 downto 3);
	s2_4(9) <= s1_5(9);
	s2_4(10) <= s1_6(10);
	s2_4(11) <= carry_2b(s1_4(10),s1_5(10));
	s2_4(12) <= carry_3b(s1_4(11),s1_5(11),s1_6(11));
	s2_4(13) <= carry_3b(s1_4(12),s1_5(12),s1_6(12));
	s2_4(14) <= carry_3b(s1_4(13),s1_5(13),s1_6(13));
	s2_4(15) <= carry_3b(s1_4(14),s1_5(14),s1_6(14));
	s2_4(16) <= carry_3b(s1_4(15),s1_5(15),s1_6(15));
	s2_4(17) <= carry_3b(s1_4(16),s1_5(16),s1_6(16));
	s2_4(18) <= carry_3b(s1_4(17),s1_5(17),s1_6(17));
	s2_4(19) <= carry_3b(s1_4(18),s1_5(18),s1_6(18));
	s2_4(20) <= carry_3b(s1_4(19),s1_5(19),s1_6(19));
	s2_4(21) <= carry_3b(s1_4(20),s1_5(20),s1_6(20));
	s2_4(22) <= carry_3b(s1_4(21),s1_5(21),s1_6(21));
	s2_4(23) <= carry_3b(s1_4(22),s1_5(22),s1_6(22));
	s2_4(24) <= carry_3b(s1_4(23),s1_5(23),s1_6(23));
	s2_4(25) <= s1_3(25);
	s2_4(29 downto 26 ) <= s1_4(29 downto 26);

	--Line 5 in 9 wires after 2nd reduction
	s2_5(8 downto 4) <= s1_5(8 downto 4);
	s2_5(9) <= s1_6(9);
	s2_5(10) <= s1_7(10);
	s2_5(11) <= sum_2b(s1_7(11),s1_8(11));
	s2_5(12) <= sum_3b(s1_7(12),s1_8(12),s1_9(12));
	s2_5(13) <= sum_3b(s1_7(13),s1_8(13),s1_9(13));
	s2_5(14) <= sum_3b(s1_7(14),s1_8(14),s1_9(14));
	s2_5(15) <= sum_3b(s1_7(15),s1_8(15),s1_9(15));
	s2_5(16) <= sum_3b(s1_7(16),s1_8(16),s1_9(16));
	s2_5(17) <= sum_3b(s1_7(17),s1_8(17),s1_9(17));
	s2_5(18) <= sum_3b(s1_7(18),s1_8(18),s1_9(18));
	s2_5(19) <= sum_3b(s1_7(19),s1_8(19),s1_9(19));
	s2_5(20) <= sum_3b(s1_7(20),s1_8(20),s1_9(20));
	s2_5(21) <= sum_3b(s1_7(21),s1_8(21),s1_9(21));
	s2_5(22) <= sum_3b(s1_7(22),s1_8(22),s1_9(22));
	s2_5(23) <= s1_7(23);
	s2_5(24) <= s1_5(24);
	s2_5(25) <= s1_4(25);
	s2_5(28 downto 26 ) <= s1_5(28 downto 26);

	--Line 6 in 9 wires after 2nd reduction
	s2_6(8 downto 5) <= s1_6(8 downto 5);
	s2_6(9) <= s1_7(9);
	s2_6(10) <= s1_8(10);
	s2_6(11) <= s1_9(11);
	s2_6(12) <= carry_2b(s1_7(11),s1_8(11));
	s2_6(13) <= carry_3b(s1_7(12),s1_8(12),s1_9(12));
	s2_6(14) <= carry_3b(s1_7(13),s1_8(13),s1_9(13));
	s2_6(15) <= carry_3b(s1_7(14),s1_8(14),s1_9(14));
	s2_6(16) <= carry_3b(s1_7(15),s1_8(15),s1_9(15));
	s2_6(17) <= carry_3b(s1_7(16),s1_8(16),s1_9(16));
	s2_6(18) <= carry_3b(s1_7(17),s1_8(17),s1_9(17));
	s2_6(19) <= carry_3b(s1_7(18),s1_8(18),s1_9(18));
	s2_6(20) <= carry_3b(s1_7(19),s1_8(19),s1_9(19));
	s2_6(21) <= carry_3b(s1_7(20),s1_8(20),s1_9(20));
	s2_6(22) <= carry_3b(s1_7(21),s1_8(21),s1_9(21));
	s2_6(23) <= carry_3b(s1_7(22),s1_8(22),s1_9(22));
	s2_6(24) <= s1_6(24);
	s2_6(25) <= s1_5(25);
	s2_6(27 downto 26 ) <= s1_6(27 downto 26);

	--Line 7 in 9 wires after 2nd reduction
	s2_7(8 downto 6) <= s1_7(8 downto 6);
	s2_7(9) <= s1_8(9);
	s2_7(10) <= s1_9(10);
	s2_7(11) <= s1_10(11);
	s2_7(12) <= sum_2b(s1_10(12),s1_11(12));
	s2_7(13) <= sum_3b(s1_10(13),s1_11(13),s1_12(13));
	s2_7(14) <= sum_3b(s1_10(14),s1_11(14),s1_12(14));
	s2_7(15) <= sum_3b(s1_10(15),s1_11(15),s1_12(15));
	s2_7(16) <= sum_3b(s1_10(16),s1_11(16),s1_12(16));
	s2_7(17) <= sum_3b(s1_10(17),s1_11(17),s1_12(17));
	s2_7(18) <= sum_3b(s1_10(18),s1_11(18),s1_12(18));
	s2_7(19) <= sum_3b(s1_10(19),s1_11(19),s1_12(19));
	s2_7(20) <= sum_3b(s1_10(20),s1_11(20),s1_12(20));
	s2_7(21) <= sum_3b(s1_10(21),s1_11(21),s1_12(21));
	s2_7(22) <= s1_10(22);
	s2_7(23) <= s1_8(23);
	s2_7(24) <= s1_7(24);
	s2_7(25) <= s1_6(25);
	s2_7(26) <= s1_7(26);

	--Line 8 in 9 wires after 2nd reduction
	s2_8(8 downto 7) <= s1_8(8 downto 7);
	s2_8(9) <= s1_9(9);
	s2_8(10) <= s1_10(10);
	s2_8(11) <= s1_11(11);
	s2_8(12) <= s1_12(12);
	s2_8(13) <= carry_2b(s1_10(12),s1_11(12));
	s2_8(14) <= carry_3b(s1_10(13),s1_11(13),s1_12(13));
	s2_8(15) <= carry_3b(s1_10(14),s1_11(14),s1_12(14));
	s2_8(16) <= carry_3b(s1_10(15),s1_11(15),s1_12(15));
	s2_8(17) <= carry_3b(s1_10(16),s1_11(16),s1_12(16));
	s2_8(18) <= carry_3b(s1_10(17),s1_11(17),s1_12(17));
	s2_8(19) <= carry_3b(s1_10(18),s1_11(18),s1_12(18));
	s2_8(20) <= carry_3b(s1_10(19),s1_11(19),s1_12(19));
	s2_8(21) <= carry_3b(s1_10(20),s1_11(20),s1_12(20));
	s2_8(22) <= carry_3b(s1_10(21),s1_11(21),s1_12(21));
	s2_8(23) <= s1_9(23);
	s2_8(24) <= s1_8(24);
	s2_8(25) <= s1_7(25);

	--Line 9 in 9 wires after 2nd reduction
	s2_9(8) <= s1_9(8);
	s2_9(9) <= s1_10(9);
	s2_9(10) <= s1_11(10);
	s2_9(11) <= s1_12(11);
	s2_9(12) <= s1_13(12);
	s2_9(21 downto 13) <= s1_13(21 downto 13);
	s2_9(22) <= s1_11(22);
	s2_9(23) <= s1_10(23);
	s2_9(24) <= s1_9(24);
	s2_9(25) <= s1_8(25);


	--Line 1 in 6 wires after 3rd reduction 
	s3_1(5 downto 0) <= s2_1(5 downto 0);
	s3_1(6 ) <= sum_2b(s2_1(6 ),s2_2(6 ));
	s3_1(7 ) <= sum_3b(s2_1(7 ),s2_2(7 ),s2_3(7));
	s3_1(8 ) <= sum_3b(s2_1(8 ),s2_2(8 ),s2_3(8));
	s3_1(9 ) <= sum_3b(s2_1(9 ),s2_2(9 ),s2_3(9));
	s3_1(10) <= sum_3b(s2_1(10),s2_2(10),s2_3(10));
	s3_1(11) <= sum_3b(s2_1(11),s2_2(11),s2_3(11));
	s3_1(12) <= sum_3b(s2_1(12),s2_2(12),s2_3(12));
	s3_1(13) <= sum_3b(s2_1(13),s2_2(13),s2_3(13));
	s3_1(14) <= sum_3b(s2_1(14),s2_2(14),s2_3(14));
	s3_1(15) <= sum_3b(s2_1(15),s2_2(15),s2_3(15));
	s3_1(16) <= sum_3b(s2_1(16),s2_2(16),s2_3(16));
	s3_1(17) <= sum_3b(s2_1(17),s2_2(17),s2_3(17));
	s3_1(18) <= sum_3b(s2_1(18),s2_2(18),s2_3(18));
	s3_1(19) <= sum_3b(s2_1(19),s2_2(19),s2_3(19));
	s3_1(20) <= sum_3b(s2_1(20),s2_2(20),s2_3(20));
	s3_1(21) <= sum_3b(s2_1(21),s2_2(21),s2_3(21));
	s3_1(22) <= sum_3b(s2_1(22),s2_2(22),s2_3(22));
	s3_1(23) <= sum_3b(s2_1(23),s2_2(23),s2_3(23));
	s3_1(24) <= sum_3b(s2_1(24),s2_2(24),s2_3(24));
	s3_1(25) <= sum_3b(s2_1(25),s2_2(25),s2_3(25));
	s3_1(26) <= sum_3b(s2_1(26),s2_2(26),s2_3(26));
	s3_1(27) <= sum_3b(s2_1(27),s2_2(27),s2_3(27));
	s3_1(32 downto 28) <= s2_1(32 downto 28);

	--Line 2 in 6 wires after 3rd reduction 
	s3_2(5 downto 1) <= s2_2(5 downto 1);
	s3_2(6) <= s2_3(6);
	s3_2(7) <= carry_2b(s2_1(6 ),s2_2(6 ));
	s3_2(8) <= carry_3b(s2_1(7 ),s2_2(7 ),s2_3(7));
	s3_2(9) <= carry_3b(s2_1(8 ),s2_2(8 ),s2_3(8));
	s3_2(10) <= carry_3b(s2_1(9 ),s2_2(9 ),s2_3(9));
	s3_2(11) <= carry_3b(s2_1(10),s2_2(10),s2_3(10));
	s3_2(12) <= carry_3b(s2_1(11),s2_2(11),s2_3(11));
	s3_2(13) <= carry_3b(s2_1(12),s2_2(12),s2_3(12));
	s3_2(14) <= carry_3b(s2_1(13),s2_2(13),s2_3(13));
	s3_2(15) <= carry_3b(s2_1(14),s2_2(14),s2_3(14));
	s3_2(16) <= carry_3b(s2_1(15),s2_2(15),s2_3(15));
	s3_2(17) <= carry_3b(s2_1(16),s2_2(16),s2_3(16));
	s3_2(18) <= carry_3b(s2_1(17),s2_2(17),s2_3(17));
	s3_2(19) <= carry_3b(s2_1(18),s2_2(18),s2_3(18));
	s3_2(20) <= carry_3b(s2_1(19),s2_2(19),s2_3(19));
	s3_2(21) <= carry_3b(s2_1(20),s2_2(20),s2_3(20));
	s3_2(22) <= carry_3b(s2_1(21),s2_2(21),s2_3(21));
	s3_2(23) <= carry_3b(s2_1(22),s2_2(22),s2_3(22));
	s3_2(24) <= carry_3b(s2_1(23),s2_2(23),s2_3(23));
	s3_2(25) <= carry_3b(s2_1(24),s2_2(24),s2_3(24));
	s3_2(26) <= carry_3b(s2_1(25),s2_2(25),s2_3(25));
	s3_2(27) <= carry_3b(s2_1(26),s2_2(26),s2_3(26));
	s3_2(28) <= carry_3b(s2_1(27),s2_2(27),s2_3(27));
	s3_2(31 downto 29) <= s2_2(31 downto 29); 


	--Line 3 in 6 wires after 3rd reduction 
	s3_3(5 downto 2) <= s2_3(5 downto 2);
	s3_3(6) <= s2_4(6);
	s3_3(7) <= sum_2b(s2_4(7),s2_5(7));
	s3_3(8) <= sum_3b(s2_4(8),s2_5(8),s2_6(8));
	s3_3(9) <= sum_3b(s2_4(9),s2_5(9),s2_6(9));
	s3_3(10) <= sum_3b(s2_4(10),s2_5(10),s2_6(10));
	s3_3(11) <= sum_3b(s2_4(11),s2_5(11),s2_6(11));
	s3_3(12) <= sum_3b(s2_4(12),s2_5(12),s2_6(12));
	s3_3(13) <= sum_3b(s2_4(13),s2_5(13),s2_6(13));
	s3_3(14) <= sum_3b(s2_4(14),s2_5(14),s2_6(14));
	s3_3(15) <= sum_3b(s2_4(15),s2_5(15),s2_6(15));
	s3_3(16) <= sum_3b(s2_4(16),s2_5(16),s2_6(16));
	s3_3(17) <= sum_3b(s2_4(17),s2_5(17),s2_6(17));
	s3_3(18) <= sum_3b(s2_4(18),s2_5(18),s2_6(18));
	s3_3(19) <= sum_3b(s2_4(19),s2_5(19),s2_6(19));
	s3_3(20) <= sum_3b(s2_4(20),s2_5(20),s2_6(20));
	s3_3(21) <= sum_3b(s2_4(21),s2_5(21),s2_6(21));
	s3_3(22) <= sum_3b(s2_4(22),s2_5(22),s2_6(22));
	s3_3(23) <= sum_3b(s2_4(23),s2_5(23),s2_6(23));
	s3_3(24) <= sum_3b(s2_4(24),s2_5(24),s2_6(24));
	s3_3(25) <= sum_3b(s2_4(25),s2_5(25),s2_6(25));
	s3_3(26) <= sum_3b(s2_4(26),s2_5(26),s2_6(26));
	s3_3(27) <= s2_4(27);
	s3_3(28) <= s2_2(28);
	s3_3(30 downto 29) <= s2_3(30 downto 29);

	--Line 4 in 6 wires after 3rd reduction 
	s3_4(5 downto 3) <= s2_4(5 downto 3);
	s3_4(6) <= s2_5(6);
	s3_4(7) <= s2_6(7);
	s3_4(8) <= carry_2b(s2_4(7),s2_5(7));
	s3_4(9) <= carry_3b(s2_4(8),s2_5(8),s2_6(8));
	s3_4(10) <= carry_3b(s2_4(9),s2_5(9),s2_6(9));
	s3_4(11) <= carry_3b(s2_4(10),s2_5(10),s2_6(10));
	s3_4(12) <= carry_3b(s2_4(11),s2_5(11),s2_6(11));
	s3_4(13) <= carry_3b(s2_4(12),s2_5(12),s2_6(12));
	s3_4(14) <= carry_3b(s2_4(13),s2_5(13),s2_6(13));
	s3_4(15) <= carry_3b(s2_4(14),s2_5(14),s2_6(14));
	s3_4(16) <= carry_3b(s2_4(15),s2_5(15),s2_6(15));
	s3_4(17) <= carry_3b(s2_4(16),s2_5(16),s2_6(16));
	s3_4(18) <= carry_3b(s2_4(17),s2_5(17),s2_6(17));
	s3_4(19) <= carry_3b(s2_4(18),s2_5(18),s2_6(18));
	s3_4(20) <= carry_3b(s2_4(19),s2_5(19),s2_6(19));
	s3_4(21) <= carry_3b(s2_4(20),s2_5(20),s2_6(20));
	s3_4(22) <= carry_3b(s2_4(21),s2_5(21),s2_6(21));
	s3_4(23) <= carry_3b(s2_4(22),s2_5(22),s2_6(22));
	s3_4(24) <= carry_3b(s2_4(23),s2_5(23),s2_6(23));
	s3_4(25) <= carry_3b(s2_4(24),s2_5(24),s2_6(24));
	s3_4(26) <= carry_3b(s2_4(25),s2_5(25),s2_6(25));
	s3_4(27) <= carry_3b(s2_4(26),s2_5(26),s2_6(26));
	s3_4(28) <= s2_3(28);
	s3_4(29) <= s2_4(29);

	--Line 5 in 6 wires after 3rd reduction 
	s3_5(5 downto 4) <= s2_5(5 downto 4);
	s3_5(6) <= s2_6(6);
	s3_5(7) <= s2_7(7);
	s3_5(8) <= sum_2b(s2_7(8),s2_8(8));
	s3_5(9) <= sum_3b(s2_7(9),s2_8(9),s2_9(9));
	s3_5(10) <= sum_3b(s2_7(10),s2_8(10),s2_9(10));
	s3_5(11) <= sum_3b(s2_7(11),s2_8(11),s2_9(11));
	s3_5(12) <= sum_3b(s2_7(12),s2_8(12),s2_9(12));
	s3_5(13) <= sum_3b(s2_7(13),s2_8(13),s2_9(13));
	s3_5(14) <= sum_3b(s2_7(14),s2_8(14),s2_9(14));
	s3_5(15) <= sum_3b(s2_7(15),s2_8(15),s2_9(15));
	s3_5(16) <= sum_3b(s2_7(16),s2_8(16),s2_9(16));
	s3_5(17) <= sum_3b(s2_7(17),s2_8(17),s2_9(17));
	s3_5(18) <= sum_3b(s2_7(18),s2_8(18),s2_9(18));
	s3_5(19) <= sum_3b(s2_7(19),s2_8(19),s2_9(19));
	s3_5(20) <= sum_3b(s2_7(20),s2_8(20),s2_9(20));
	s3_5(21) <= sum_3b(s2_7(21),s2_8(21),s2_9(21));
	s3_5(22) <= sum_3b(s2_7(22),s2_8(22),s2_9(22));
	s3_5(23) <= sum_3b(s2_7(23),s2_8(23),s2_9(23));
	s3_5(24) <= sum_3b(s2_7(24),s2_8(24),s2_9(24));
	s3_5(25) <= sum_3b(s2_7(25),s2_8(25),s2_9(25));
	s3_5(26) <= s2_7(26);
	s3_5(27) <= s2_5(27);
	s3_5(28) <= s2_4(28);

	--Line 6 in 6 wires after 3rd reduction 
	s3_6(5) <= s2_6(5);
	s3_6(6) <= s2_7(6);
	s3_6(7) <= s2_8(7);
	s3_6(8) <= s2_9(8);
	s3_6(9) <= carry_2b(s2_7(8),s2_8(8));
	s3_6(10) <= carry_3b(s2_7(9),s2_8(9),s2_9(9));
	s3_6(11) <= carry_3b(s2_7(10),s2_8(10),s2_9(10));
	s3_6(12) <= carry_3b(s2_7(11),s2_8(11),s2_9(11));
	s3_6(13) <= carry_3b(s2_7(12),s2_8(12),s2_9(12));
	s3_6(14) <= carry_3b(s2_7(13),s2_8(13),s2_9(13));
	s3_6(15) <= carry_3b(s2_7(14),s2_8(14),s2_9(14));
	s3_6(16) <= carry_3b(s2_7(15),s2_8(15),s2_9(15));
	s3_6(17) <= carry_3b(s2_7(16),s2_8(16),s2_9(16));
	s3_6(18) <= carry_3b(s2_7(17),s2_8(17),s2_9(17));
	s3_6(19) <= carry_3b(s2_7(18),s2_8(18),s2_9(18));
	s3_6(20) <= carry_3b(s2_7(19),s2_8(19),s2_9(19));
	s3_6(21) <= carry_3b(s2_7(20),s2_8(20),s2_9(20));
	s3_6(22) <= carry_3b(s2_7(21),s2_8(21),s2_9(21));
	s3_6(23) <= carry_3b(s2_7(22),s2_8(22),s2_9(22));
	s3_6(24) <= carry_3b(s2_7(23),s2_8(23),s2_9(23));
	s3_6(25) <= carry_3b(s2_7(24),s2_8(24),s2_9(24));
	s3_6(26) <= carry_3b(s2_7(25),s2_8(25),s2_9(25));
	s3_6(27) <= s2_6(27);
	s3_6(28) <= s2_5(28);


	--Line 1 in 4 wires after 4th reduction 
	s4_1(3 downto 0) <= s3_1(3 downto 0);
	s4_1(4) <= sum_2b(s3_1(4),s3_2(4));
	s4_1(5 ) <= sum_3b(s3_1(5),s3_2(5),s3_3(5));
	s4_1(6 ) <= sum_3b(s3_1(6),s3_2(6),s3_3(6));
	s4_1(7 ) <= sum_3b(s3_1(7),s3_2(7),s3_3(7));
	s4_1(8 ) <= sum_3b(s3_1(8),s3_2(8),s3_3(8));
	s4_1(9 ) <= sum_3b(s3_1(9),s3_2(9),s3_3(9));
	s4_1(10) <= sum_3b(s3_1(10),s3_2(10),s3_3(10));
	s4_1(11) <= sum_3b(s3_1(11),s3_2(11),s3_3(11));
	s4_1(12) <= sum_3b(s3_1(12),s3_2(12),s3_3(12));
	s4_1(13) <= sum_3b(s3_1(13),s3_2(13),s3_3(13));
	s4_1(14) <= sum_3b(s3_1(14),s3_2(14),s3_3(14));
	s4_1(15) <= sum_3b(s3_1(15),s3_2(15),s3_3(15));
	s4_1(16) <= sum_3b(s3_1(16),s3_2(16),s3_3(16));
	s4_1(17) <= sum_3b(s3_1(17),s3_2(17),s3_3(17));
	s4_1(18) <= sum_3b(s3_1(18),s3_2(18),s3_3(18));
	s4_1(19) <= sum_3b(s3_1(19),s3_2(19),s3_3(19));
	s4_1(20) <= sum_3b(s3_1(20),s3_2(20),s3_3(20));
	s4_1(21) <= sum_3b(s3_1(21),s3_2(21),s3_3(21));
	s4_1(22) <= sum_3b(s3_1(22),s3_2(22),s3_3(22));
	s4_1(23) <= sum_3b(s3_1(23),s3_2(23),s3_3(23));
	s4_1(24) <= sum_3b(s3_1(24),s3_2(24),s3_3(24));
	s4_1(25) <= sum_3b(s3_1(25),s3_2(25),s3_3(25));
	s4_1(26) <= sum_3b(s3_1(26),s3_2(26),s3_3(26));
	s4_1(27) <= sum_3b(s3_1(27),s3_2(27),s3_3(27));
	s4_1(28) <= sum_3b(s3_1(28),s3_2(28),s3_3(28));
	s4_1(29) <= sum_3b(s3_1(29),s3_2(29),s3_3(29));
	s4_1(32 downto 30) <= s3_1(32 downto 30);

	--Line 2 in 4 wires after 4th reduction 
	s4_2(3 downto 1) <= s3_2(3 downto 1);
	s4_2(4) <= s3_3(4);
	s4_2(5) <= carry_2b(s3_1(4),s3_2(4));
	s4_2(6 ) <= carry_3b(s3_1(5),s3_2(5),s3_3(5));
	s4_2(7 ) <= carry_3b(s3_1(6),s3_2(6),s3_3(6));
	s4_2(8 ) <= carry_3b(s3_1(7),s3_2(7),s3_3(7));
	s4_2(9 ) <= carry_3b(s3_1(8),s3_2(8),s3_3(8));
	s4_2(10) <= carry_3b(s3_1(9),s3_2(9),s3_3(9));
	s4_2(11) <= carry_3b(s3_1(10),s3_2(10),s3_3(10));
	s4_2(12) <= carry_3b(s3_1(11),s3_2(11),s3_3(11));
	s4_2(13) <= carry_3b(s3_1(12),s3_2(12),s3_3(12));
	s4_2(14) <= carry_3b(s3_1(13),s3_2(13),s3_3(13));
	s4_2(15) <= carry_3b(s3_1(14),s3_2(14),s3_3(14));
	s4_2(16) <= carry_3b(s3_1(15),s3_2(15),s3_3(15));
	s4_2(17) <= carry_3b(s3_1(16),s3_2(16),s3_3(16));
	s4_2(18) <= carry_3b(s3_1(17),s3_2(17),s3_3(17));
	s4_2(19) <= carry_3b(s3_1(18),s3_2(18),s3_3(18));
	s4_2(20) <= carry_3b(s3_1(19),s3_2(19),s3_3(19));
	s4_2(21) <= carry_3b(s3_1(20),s3_2(20),s3_3(20));
	s4_2(22) <= carry_3b(s3_1(21),s3_2(21),s3_3(21));
	s4_2(23) <= carry_3b(s3_1(22),s3_2(22),s3_3(22));
	s4_2(24) <= carry_3b(s3_1(23),s3_2(23),s3_3(23));
	s4_2(25) <= carry_3b(s3_1(24),s3_2(24),s3_3(24));
	s4_2(26) <= carry_3b(s3_1(25),s3_2(25),s3_3(25));
	s4_2(27) <= carry_3b(s3_1(26),s3_2(26),s3_3(26));
	s4_2(28) <= carry_3b(s3_1(27),s3_2(27),s3_3(27));
	s4_2(29) <= carry_3b(s3_1(28),s3_2(28),s3_3(28));
	s4_2(30) <= carry_3b(s3_1(29),s3_2(29),s3_3(29));
	s4_2(31) <= s3_2(31);

	--Line 3 in 4 wires after 4th reduction 
	s4_3(3 downto 2) <= s3_3(3 downto 2);
	s4_3(4) <= s3_4(4);
	s4_3(5) <= sum_2b(s3_4(5),s3_5(5));
	s4_3(6 ) <= sum_3b(s3_4(6 ),s3_5(6 ),s3_6(6 ));
	s4_3(7 ) <= sum_3b(s3_4(7 ),s3_5(7 ),s3_6(7 ));
	s4_3(8 ) <= sum_3b(s3_4(8 ),s3_5(8 ),s3_6(8 ));
	s4_3(9 ) <= sum_3b(s3_4(9 ),s3_5(9 ),s3_6(9 ));
	s4_3(10) <= sum_3b(s3_4(10),s3_5(10),s3_6(10));
	s4_3(11) <= sum_3b(s3_4(11),s3_5(11),s3_6(11));
	s4_3(12) <= sum_3b(s3_4(12),s3_5(12),s3_6(12));
	s4_3(13) <= sum_3b(s3_4(13),s3_5(13),s3_6(13));
	s4_3(14) <= sum_3b(s3_4(14),s3_5(14),s3_6(14));
	s4_3(15) <= sum_3b(s3_4(15),s3_5(15),s3_6(15));
	s4_3(16) <= sum_3b(s3_4(16),s3_5(16),s3_6(16));
	s4_3(17) <= sum_3b(s3_4(17),s3_5(17),s3_6(17));
	s4_3(18) <= sum_3b(s3_4(18),s3_5(18),s3_6(18));
	s4_3(19) <= sum_3b(s3_4(19),s3_5(19),s3_6(19));
	s4_3(20) <= sum_3b(s3_4(20),s3_5(20),s3_6(20));
	s4_3(21) <= sum_3b(s3_4(21),s3_5(21),s3_6(21));
	s4_3(22) <= sum_3b(s3_4(22),s3_5(22),s3_6(22));
	s4_3(23) <= sum_3b(s3_4(23),s3_5(23),s3_6(23));
	s4_3(24) <= sum_3b(s3_4(24),s3_5(24),s3_6(24));
	s4_3(25) <= sum_3b(s3_4(25),s3_5(25),s3_6(25));
	s4_3(26) <= sum_3b(s3_4(26),s3_5(26),s3_6(26));
	s4_3(27) <= sum_3b(s3_4(27),s3_5(27),s3_6(27));
	s4_3(28) <= sum_3b(s3_4(28),s3_5(28),s3_6(28));
	s4_3(29) <= s3_4(29);
	s4_3(30) <= s3_2(30);

	--Line 4 in 4 wires after 4th reduction 
	s4_4(3) <= s3_4(3);
	s4_4(4) <= s3_5(4);
	s4_4(5) <= s3_6(5);
	s4_4(6) <= carry_2b(s3_4(5),s3_5(5));
	s4_4(7) <= carry_3b(s3_4(6 ),s3_5(6 ),s3_6(6 ));
	s4_4(8) <= carry_3b(s3_4(7 ),s3_5(7 ),s3_6(7 ));
	s4_4(9) <= carry_3b(s3_4(8 ),s3_5(8 ),s3_6(8 ));
	s4_4(10) <= carry_3b(s3_4(9 ),s3_5(9 ),s3_6(9 ));
	s4_4(11) <= carry_3b(s3_4(10),s3_5(10),s3_6(10));
	s4_4(12) <= carry_3b(s3_4(11),s3_5(11),s3_6(11));
	s4_4(13) <= carry_3b(s3_4(12),s3_5(12),s3_6(12));
	s4_4(14) <= carry_3b(s3_4(13),s3_5(13),s3_6(13));
	s4_4(15) <= carry_3b(s3_4(14),s3_5(14),s3_6(14));
	s4_4(16) <= carry_3b(s3_4(15),s3_5(15),s3_6(15));
	s4_4(17) <= carry_3b(s3_4(16),s3_5(16),s3_6(16));
	s4_4(18) <= carry_3b(s3_4(17),s3_5(17),s3_6(17));
	s4_4(19) <= carry_3b(s3_4(18),s3_5(18),s3_6(18));
	s4_4(20) <= carry_3b(s3_4(19),s3_5(19),s3_6(19));
	s4_4(21) <= carry_3b(s3_4(20),s3_5(20),s3_6(20));
	s4_4(22) <= carry_3b(s3_4(21),s3_5(21),s3_6(21));
	s4_4(23) <= carry_3b(s3_4(22),s3_5(22),s3_6(22));
	s4_4(24) <= carry_3b(s3_4(23),s3_5(23),s3_6(23));
	s4_4(25) <= carry_3b(s3_4(24),s3_5(24),s3_6(24));
	s4_4(26) <= carry_3b(s3_4(25),s3_5(25),s3_6(25));
	s4_4(27) <= carry_3b(s3_4(26),s3_5(26),s3_6(26));
	s4_4(28) <= carry_3b(s3_4(27),s3_5(27),s3_6(27));
	s4_4(29) <= carry_3b(s3_4(28),s3_5(28),s3_6(28));
	s4_4(30) <= s3_3(30);

	--Line 1 in 3 wires after 5th reduction
	s5_1(2 downto 0) <= s4_1(2 downto 0);
	s5_1(3) <= sum_2b(s4_1(3),s4_2(3));
	s5_1(4) <= sum_3b(s4_1(4),s4_2(4),s4_3(4));
	s5_1(5) <= sum_3b(s4_1(5),s4_2(5),s4_3(5));
	s5_1(6) <= sum_3b(s4_1(6),s4_2(6),s4_3(6));
	s5_1(7) <= sum_3b(s4_1(7),s4_2(7),s4_3(7));
	s5_1(8) <= sum_3b(s4_1(8),s4_2(8),s4_3(8));
	s5_1(9) <= sum_3b(s4_1(9),s4_2(9),s4_3(9));
	s5_1(10) <= sum_3b(s4_1(10),s4_2(10),s4_3(10));
	s5_1(11) <= sum_3b(s4_1(11),s4_2(11),s4_3(11));
	s5_1(12) <= sum_3b(s4_1(12),s4_2(12),s4_3(12));
	s5_1(13) <= sum_3b(s4_1(13),s4_2(13),s4_3(13));
	s5_1(14) <= sum_3b(s4_1(14),s4_2(14),s4_3(14));
	s5_1(15) <= sum_3b(s4_1(15),s4_2(15),s4_3(15));
	s5_1(16) <= sum_3b(s4_1(16),s4_2(16),s4_3(16));
	s5_1(17) <= sum_3b(s4_1(17),s4_2(17),s4_3(17));
	s5_1(18) <= sum_3b(s4_1(18),s4_2(18),s4_3(18));
	s5_1(19) <= sum_3b(s4_1(19),s4_2(19),s4_3(19));
	s5_1(20) <= sum_3b(s4_1(20),s4_2(20),s4_3(20));
	s5_1(21) <= sum_3b(s4_1(21),s4_2(21),s4_3(21));
	s5_1(22) <= sum_3b(s4_1(22),s4_2(22),s4_3(22));
	s5_1(23) <= sum_3b(s4_1(23),s4_2(23),s4_3(23));
	s5_1(24) <= sum_3b(s4_1(24),s4_2(24),s4_3(24));
	s5_1(25) <= sum_3b(s4_1(25),s4_2(25),s4_3(25));
	s5_1(26) <= sum_3b(s4_1(26),s4_2(26),s4_3(26));
	s5_1(27) <= sum_3b(s4_1(27),s4_2(27),s4_3(27));
	s5_1(28) <= sum_3b(s4_1(28),s4_2(28),s4_3(28));
	s5_1(29) <= sum_3b(s4_1(29),s4_2(29),s4_3(29));
	s5_1(30) <= sum_3b(s4_1(30),s4_2(30),s4_3(30));
	s5_1(31) <= s4_1(31);
	s5_1(32) <= s4_1(32);

	--Line 2 in 3 wires after 5th reduction
	s5_2(2 downto 1) <= s4_2(2 downto 1);
	s5_2(3) <= s4_3(3);
	s5_2(4) <= carry_2b(s4_1(3),s4_2(3));
	s5_2(5) <= carry_3b(s4_1(4),s4_2(4),s4_3(4));
	s5_2(6) <= carry_3b(s4_1(5),s4_2(5),s4_3(5));
	s5_2(7) <= carry_3b(s4_1(6),s4_2(6),s4_3(6));
	s5_2(8) <= carry_3b(s4_1(7),s4_2(7),s4_3(7));
	s5_2(9) <= carry_3b(s4_1(8),s4_2(8),s4_3(8));
	s5_2(10) <= carry_3b(s4_1(9),s4_2(9),s4_3(9));
	s5_2(11) <= carry_3b(s4_1(10),s4_2(10),s4_3(10));
	s5_2(12) <= carry_3b(s4_1(11),s4_2(11),s4_3(11));
	s5_2(13) <= carry_3b(s4_1(12),s4_2(12),s4_3(12));
	s5_2(14) <= carry_3b(s4_1(13),s4_2(13),s4_3(13));
	s5_2(15) <= carry_3b(s4_1(14),s4_2(14),s4_3(14));
	s5_2(16) <= carry_3b(s4_1(15),s4_2(15),s4_3(15));
	s5_2(17) <= carry_3b(s4_1(16),s4_2(16),s4_3(16));
	s5_2(18) <= carry_3b(s4_1(17),s4_2(17),s4_3(17));
	s5_2(19) <= carry_3b(s4_1(18),s4_2(18),s4_3(18));
	s5_2(20) <= carry_3b(s4_1(19),s4_2(19),s4_3(19));
	s5_2(21) <= carry_3b(s4_1(20),s4_2(20),s4_3(20));
	s5_2(22) <= carry_3b(s4_1(21),s4_2(21),s4_3(21));
	s5_2(23) <= carry_3b(s4_1(22),s4_2(22),s4_3(22));
	s5_2(24) <= carry_3b(s4_1(23),s4_2(23),s4_3(23));
	s5_2(25) <= carry_3b(s4_1(24),s4_2(24),s4_3(24));
	s5_2(26) <= carry_3b(s4_1(25),s4_2(25),s4_3(25));
	s5_2(27) <= carry_3b(s4_1(26),s4_2(26),s4_3(26));
	s5_2(28) <= carry_3b(s4_1(27),s4_2(27),s4_3(27));
	s5_2(29) <= carry_3b(s4_1(28),s4_2(28),s4_3(28));
	s5_2(30) <= carry_3b(s4_1(29),s4_2(29),s4_3(29));
	s5_2(31) <= carry_3b(s4_1(30),s4_2(30),s4_3(30));
	
	--Line 3 in 3 wires after 5th reduction
	s5_3(2) <= s4_3(2);
	s5_3(30 downto 3) <= s4_4(30 downto 3);
	s5_3(31) <= s4_2(31);

	--Line 1 in 2 wires after 6th reduction 
	s6_1(1 downto 0) <= s5_1(1 downto 0);
	s6_1(2) <= sum_2b(s5_1(2),s5_2(2));
	s6_1(3) <= sum_3b(s5_1(3),s5_2(3),s5_3(3));
	s6_1(4) <= sum_3b(s5_1(4),s5_2(4),s5_3(4));
	s6_1(5) <= sum_3b(s5_1(5),s5_2(5),s5_3(5));
	s6_1(6) <= sum_3b(s5_1(6),s5_2(6),s5_3(6));
	s6_1(7) <= sum_3b(s5_1(7),s5_2(7),s5_3(7));
	s6_1(8) <= sum_3b(s5_1(8),s5_2(8),s5_3(8));
	s6_1(9) <= sum_3b(s5_1(9),s5_2(9),s5_3(9));
	s6_1(10) <= sum_3b(s5_1(10),s5_2(10),s5_3(10));
	s6_1(11) <= sum_3b(s5_1(11),s5_2(11),s5_3(11));
	s6_1(12) <= sum_3b(s5_1(12),s5_2(12),s5_3(12));
	s6_1(13) <= sum_3b(s5_1(13),s5_2(13),s5_3(13));
	s6_1(14) <= sum_3b(s5_1(14),s5_2(14),s5_3(14));
	s6_1(15) <= sum_3b(s5_1(15),s5_2(15),s5_3(15));
	s6_1(16) <= sum_3b(s5_1(16),s5_2(16),s5_3(16));
	s6_1(17) <= sum_3b(s5_1(17),s5_2(17),s5_3(17));
	s6_1(18) <= sum_3b(s5_1(18),s5_2(18),s5_3(18));
	s6_1(19) <= sum_3b(s5_1(19),s5_2(19),s5_3(19));
	s6_1(20) <= sum_3b(s5_1(20),s5_2(20),s5_3(20));
	s6_1(21) <= sum_3b(s5_1(21),s5_2(21),s5_3(21));
	s6_1(22) <= sum_3b(s5_1(22),s5_2(22),s5_3(22));
	s6_1(23) <= sum_3b(s5_1(23),s5_2(23),s5_3(23));
	s6_1(24) <= sum_3b(s5_1(24),s5_2(24),s5_3(24));
	s6_1(25) <= sum_3b(s5_1(25),s5_2(25),s5_3(25));
	s6_1(26) <= sum_3b(s5_1(26),s5_2(26),s5_3(26));
	s6_1(27) <= sum_3b(s5_1(27),s5_2(27),s5_3(27));
	s6_1(28) <= sum_3b(s5_1(28),s5_2(28),s5_3(28));
	s6_1(29) <= sum_3b(s5_1(29),s5_2(29),s5_3(29));
	s6_1(30) <= sum_3b(s5_1(30),s5_2(30),s5_3(30));
	s6_1(31) <= sum_3b(s5_1(31),s5_2(31),s5_3(31));
	s6_1(32) <= s5_1(32);

	--Line 2 in 2 wires after 6th reduction 
	S6_2(0) <= '0';
	s6_2(1) <= s5_2(1);
	s6_2(2) <= s5_3(2);
	s6_2(3) <= carry_2b(s5_1(2),s5_2(2));
	s6_2(4) <= carry_3b(s5_1(3),s5_2(3),s5_3(3));
	s6_2(5) <= carry_3b(s5_1(4),s5_2(4),s5_3(4));
	s6_2(6) <= carry_3b(s5_1(5),s5_2(5),s5_3(5));
	s6_2(7) <= carry_3b(s5_1(6),s5_2(6),s5_3(6));
	s6_2(8) <= carry_3b(s5_1(7),s5_2(7),s5_3(7));
	s6_2(9) <= carry_3b(s5_1(8),s5_2(8),s5_3(8));
	s6_2(10) <= carry_3b(s5_1(9),s5_2(9),s5_3(9));
	s6_2(11) <= carry_3b(s5_1(10),s5_2(10),s5_3(10));
	s6_2(12) <= carry_3b(s5_1(11),s5_2(11),s5_3(11));
	s6_2(13) <= carry_3b(s5_1(12),s5_2(12),s5_3(12));
	s6_2(14) <= carry_3b(s5_1(13),s5_2(13),s5_3(13));
	s6_2(15) <= carry_3b(s5_1(14),s5_2(14),s5_3(14));
	s6_2(16) <= carry_3b(s5_1(15),s5_2(15),s5_3(15));
	s6_2(17) <= carry_3b(s5_1(16),s5_2(16),s5_3(16));
	s6_2(18) <= carry_3b(s5_1(17),s5_2(17),s5_3(17));
	s6_2(19) <= carry_3b(s5_1(18),s5_2(18),s5_3(18));
	s6_2(20) <= carry_3b(s5_1(19),s5_2(19),s5_3(19));
	s6_2(21) <= carry_3b(s5_1(20),s5_2(20),s5_3(20));
	s6_2(22) <= carry_3b(s5_1(21),s5_2(21),s5_3(21));
	s6_2(23) <= carry_3b(s5_1(22),s5_2(22),s5_3(22));
	s6_2(24) <= carry_3b(s5_1(23),s5_2(23),s5_3(23));
	s6_2(25) <= carry_3b(s5_1(24),s5_2(24),s5_3(24));
	s6_2(26) <= carry_3b(s5_1(25),s5_2(25),s5_3(25));
	s6_2(27) <= carry_3b(s5_1(26),s5_2(26),s5_3(26));
	s6_2(28) <= carry_3b(s5_1(27),s5_2(27),s5_3(27));
	s6_2(29) <= carry_3b(s5_1(28),s5_2(28),s5_3(28));
	s6_2(30) <= carry_3b(s5_1(29),s5_2(29),s5_3(29));
	s6_2(31) <= carry_3b(s5_1(30),s5_2(30),s5_3(30));
	s6_2(32) <= carry_3b(s5_1(31),s5_2(31),s5_3(31));

	--Final Addition
	p(32 downto 0) <= std_logic_vector(unsigned(s6_1(32 downto 0)) + unsigned(s6_2(32 downto 0)));
	p(33) <= a(16) xor b(16);
end architecture;
